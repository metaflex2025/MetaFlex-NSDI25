-- find first  library ieee;use ieee.std_logic_1164.all;use ieee.numeric_std.all;use ieee.std_logic_misc.all;use IEEE.math_real.all;entity tb_find_earliest_non_empty_fifo_1k isend tb_find_earliest_non_empty_fifo_1k;architecture test_bench of tb_find_earliest_non_empty_fifo_1k isconstant g_L2_FIFO_NUM      : integer := 10;constant g_FIFO_NUM         : integer := 2**g_L2_FIFO_NUM;constant g_L2_LEAF_FIFO_NUM : integer := 5;constant g_LEAF_FIFO_NUM    : integer := 2**g_L2_LEAF_FIFO_NUM;component find_earliest_non_empty_fifo_1k is  generic (    g_L2_FIFO_NUM       : integer;     -- log2 of number of FIFOs    g_FIFO_NUM          : integer      -- Number of FIFOs  );  port (    rst                              : in  std_logic;    clk                              : in  std_logic;    find_earliest_non_empty_fifo_cmd : in  std_logic;    current_fifo_index               : in  unsigned(g_L2_FIFO_NUM - 1 downto 0);    empty                            : in  std_logic_vector(g_FIFO_NUM-1 downto 0);    find_earliest_non_empty_fifo_rsp : out std_logic;    earliest_fifo_index              : out unsigned(g_L2_FIFO_NUM - 1 downto 0);    all_fifos_empty                  : out std_logic  );end component find_earliest_non_empty_fifo_1k;signal rst : std_logic := '0';signal clk : std_logic := '0';signal find_earliest_non_empty_fifo_cmd : std_logic := '0';signal current_fifo_index: unsigned(g_L2_FIFO_NUM - 1 downto 0) := (others => '0');signal empty : std_logic_vector(g_FIFO_NUM - 1 downto 0) := (others => '1');signal find_earliest_non_empty_fifo_rsp : std_logic;signal earliest_fifo_index : unsigned(g_L2_FIFO_NUM - 1 downto 0);signal all_fifos_empty : std_logic;beginprocessbegin    wait for 2 ns;    rst <= '1';    wait for 2 ns;    rst <= '0';    wait;end process;processbegin    for t in 0 to 50    loop        clk <= not clk;        wait for 1 ns;    end loop;    wait;end process;processbegin    wait for 0.1 ns;    wait for 4 ns;        -- Earliest FF = 1    find_earliest_non_empty_fifo_cmd <= '1';    empty <= (1023 downto 2 => '1') & '0' & '1';    wait for 2 ns;    find_earliest_non_empty_fifo_cmd <= '0';    wait for 4 ns;        -- Earliest FF = 35    find_earliest_non_empty_fifo_cmd <= '1';    empty <= (1023 downto 36 => '1') & '0' & (34 downto 0 => '1');    wait for 2 ns;    find_earliest_non_empty_fifo_cmd <= '0';    wait for 4 ns;        -- Earliest FF = 101    current_fifo_index <= to_unsigned(31, g_L2_FIFO_NUM);        find_earliest_non_empty_fifo_cmd <= '1';    empty <= (1023 downto 102 => '1') & '0' & (100 downto 2 => '1') & '0' & '1';    wait for 2 ns;    find_earliest_non_empty_fifo_cmd <= '0';    wait for 4 ns;        -- Earliest FF = 1       current_fifo_index <= to_unsigned(102, g_L2_FIFO_NUM);        find_earliest_non_empty_fifo_cmd <= '1';    empty <= (1023 downto 102 => '1') & '0' & (100 downto 2 => '1') & '0' & '1';    wait for 2 ns;    find_earliest_non_empty_fifo_cmd <= '0';    wait for 4 ns;        wait;end process;ff_1k_ii: find_earliest_non_empty_fifo_1k  generic map (    g_L2_FIFO_NUM      => g_L2_FIFO_NUM,     -- log2 of number of FIFOs    g_FIFO_NUM         => g_FIFO_NUM         -- Number of FIFOs  )  port map (    rst                              => rst,    clk                              => clk,    find_earliest_non_empty_fifo_cmd => find_earliest_non_empty_fifo_cmd,    current_fifo_index               => current_fifo_index,    empty                            => empty,    find_earliest_non_empty_fifo_rsp => find_earliest_non_empty_fifo_rsp,    earliest_fifo_index              => earliest_fifo_index,    all_fifos_empty                  => all_fifos_empty  );end test_bench; 